library verilog;
use verilog.vl_types.all;
entity VectorProcessor_tb is
end VectorProcessor_tb;
